-- Top level disign of rsa crpyto core


library ieee;
use ieee.std_logic_1164.all;


entity RSACore is
	port (
		Clk 		: in std_logic;
		Resetn 		: in std_logic);
		


end RSACCore;
